module rtl();
endmodule
