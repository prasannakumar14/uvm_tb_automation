package pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "xtn.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "sequencer.sv"
  `include "agent.sv"
  `include "sequence.sv"

  `include "env.sv"
  `include "test.sv"
endpackage
